`timescale 1ns / 1ps
`default_nettype none

module com_tb;
    //make logics for inputs and outputs!
    stereo_match uut();

    always begin
    end

    initial begin
        
    end

endmodule

`default_nettype wire