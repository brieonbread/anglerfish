/***********************************************************************
 * An RTL model of a 10-to-4 Priority BCD Encoder.
 *
 * SystemVerilog Training Workshop.
 *
 * Copyright by Sutherland HDL, Inc.
 * Tualatin, Oregon, USA.
 * www.sutherland-hdl.com
 * All rights reserved.
 **********************************************************************/

module bcd_encoder (
  input  logic [9:1] decimal_in,
  output logic [3:0] bcd_out
);
  timeunit 1ns; timeprecision 1ns;

  always_comb begin
  // ADD 10-line to 4-line PRIORITY BCD ENCODER FUNCTIONALITY

  end
endmodule
